module and1(o, x, y);
output o;
input x, y;

and x1(o, x, y)

endmodule